module stable_input (clk, reset, in, out);
	input logic clk, reset, in;
	output logic out;
	
endmodule
